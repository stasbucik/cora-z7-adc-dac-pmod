----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/31/2025 02:26:07 PM
-- Design Name: 
-- Module Name: Axi4InterfaceTb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

use std.env.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

use IEEE.math_real."ceil";
use IEEE.math_real."log2";

use work.BramPkg.all;
use work.BramBufferPkg.all;
use work.Axi4Pkg.all;

use std.textio.all;

entity Axi4InterfaceTb is
--  Port ( );
end Axi4InterfaceTb;

architecture Behavioral of Axi4InterfaceTb is

	constant CLK_PERIOD_C        : time    := 10 ns;
	constant TB_AXI_DATA_WIDTH_C : natural := 32;
	constant TB_AXI_ADDR_WIDTH_C : natural := 32;

	constant TB_NUM_ADDRESSES_C     : natural := 8;
	constant TB_PACKING_C           : natural := 2;
	constant TB_SAMPLE_DATA_WIDTH_C : natural := 12;
	constant TB_DATA_WIDTH_C        : natural := TB_PACKING_C * TB_SAMPLE_DATA_WIDTH_C;
	constant TB_BYTE_WIDTH_C        : natural := TB_DATA_WIDTH_C;
	constant TB_LATENCY_C           : natural := 3;
	constant TB_MEMORY_SIZE_C       : natural := TB_NUM_ADDRESSES_C * TB_DATA_WIDTH_C;
	constant TB_ADDR_WIDTH_C        : natural := natural(ceil(log2(real(TB_NUM_ADDRESSES_C))));
	constant TB_MAX_LENGTH_C        : natural := 256;
	constant TB_LENGTH_WIDTH_C      : natural := natural(ceil(log2(real(TB_MAX_LENGTH_C))));

	-- UUT signals
	signal clk_i : STD_LOGIC;
	signal rst_i : STD_LOGIC;
	signal axiReadSrc_i : Axi4ReadSource;
	signal axiReadDst_o : Axi4ReadDestination;
	signal readStart_o  : STD_LOGIC;
	signal address_o    : STD_LOGIC_VECTOR(TB_ADDR_WIDTH_C-1 downto 0);
	signal length_o     : STD_LOGIC_VECTOR(TB_LENGTH_WIDTH_C-1 downto 0);
	signal readDone_i   : STD_LOGIC;
	signal counter_i    : unsigned(TB_LENGTH_WIDTH_C-1 downto 0);
	signal buffer_i     : TmpBufferArray(TB_MAX_LENGTH_C-1 downto 0)(TB_DATA_WIDTH_C-1 downto 0);

	constant AXI_READ_SRC_INIT_C : axiReadSrc_i'subtype := (
			ARID     => (others => '0'),
			ARADDR   => (others => '0'),
			ARLEN    => (others => '0'),
			ARSIZE   => (others => '0'),
			ARBURST  => (others => '0'),
			ARLOCK   => (others => '0'),
			ARCACHE  => (others => '0'),
			ARPROT   => (others => '0'),
			ARQOS    => (others => '0'),
			ARREGION => (others => '0'),
			ARUSER   => (others => '0'),
			ARVALID  => '0',
			RREADY   => '0'
		);

begin

	clock : process
	begin
		clk_i <= '1';
		wait for CLK_PERIOD_C/2;
		clk_i <= '0';
		wait for CLK_PERIOD_C/2;
	end process;

	-- UUT
	Axi4Interface_1 : entity work.Axi4Interface
		generic map (
			PACKING_G           => TB_PACKING_C,
			SAMPLE_DATA_WIDTH_G => TB_SAMPLE_DATA_WIDTH_C,
			DATA_WIDTH_G        => TB_DATA_WIDTH_C,
			MAX_LENGTH_G        => TB_MAX_LENGTH_C,
			LENGTH_WIDTH_G      => TB_LENGTH_WIDTH_C,
			ADDR_WIDTH_G        => TB_ADDR_WIDTH_C
		)
		port map (
			clk_i        => clk_i,
			rst_i        => rst_i,
			axiReadSrc_i => axiReadSrc_i,
			axiReadDst_o => axiReadDst_o,
			readStart_o  => readStart_o,
			address_o    => address_o,
			length_o     => length_o,
			readDone_i   => readDone_i,
			counter_i    => counter_i,
			buffer_i     => buffer_i
		);

	stimulus : process
	begin
		rst_i <= '1';
		-- initialize signals
		axiReadSrc_i <= AXI_READ_SRC_INIT_C;

		readDone_i <= '0';
		counter_i  <= (others => '0');
		buffer_i   <= (others => (others => '0'));

		wait for CLK_PERIOD_C*3;
		rst_i <= '0';
		------------------------------------------------------------------------
		-- reset done
		------------------------------------------------------------------------
		wait for CLK_PERIOD_C*5;

		-- axi ready immediately, wait for data, read 1
		axiReadSrc_i.araddr  <= STD_LOGIC_VECTOR(to_unsigned(0, axiReadSrc_i.araddr'length));
		axiReadSrc_i.arlen   <= STD_LOGIC_VECTOR(to_unsigned(1-1, axiReadSrc_i.arlen'length));
		axiReadSrc_i.arsize  <= "101";
		axiReadSrc_i.arburst <= "01";
		axiReadSrc_i.arvalid <= '1';
		axiReadSrc_i.rready  <= '1';
		wait for CLK_PERIOD_C;
		axiReadSrc_i.arvalid <= '0';

		wait for CLK_PERIOD_C * 10;
		counter_i   <= to_unsigned(1, counter_i'length);
		readDone_i  <= '1';
		buffer_i(0) <= x"badb17";

		wait until axiReadDst_o.rvalid = '1';
		wait for CLK_PERIOD_C;
		readDone_i           <= '0';
		counter_i            <= (others => '0');
		buffer_i             <= (others => (others => '0'));
		axiReadSrc_i.araddr  <= (others => '0');
		axiReadSrc_i.arlen   <= (others => '0');
		axiReadSrc_i.arsize  <= "000";
		axiReadSrc_i.arburst <= "00";
		axiReadSrc_i.arvalid <= '0';
		axiReadSrc_i.rready  <= '0';
		wait for CLK_PERIOD_C * 5;



		-- axi not ready immediately, data is availible immediately, read 1
		axiReadSrc_i.araddr  <= STD_LOGIC_VECTOR(to_unsigned(0, axiReadSrc_i.araddr'length));
		axiReadSrc_i.arlen   <= STD_LOGIC_VECTOR(to_unsigned(1-1, axiReadSrc_i.arlen'length));
		axiReadSrc_i.arsize  <= "101";
		axiReadSrc_i.arburst <= "01";
		axiReadSrc_i.arvalid <= '1';
		wait for CLK_PERIOD_C;
		axiReadSrc_i.arvalid <= '0';

		wait for CLK_PERIOD_C * 2;
		counter_i   <= to_unsigned(1, counter_i'length);
		readDone_i  <= '1';
		buffer_i(0) <= x"badb17";

		wait for CLK_PERIOD_C * 10;
		axiReadSrc_i.rready <= '1';

		report "rvalid: " & STD_LOGIC'image(axiReadDst_o.rvalid);
		--wait until axiReadDst_o.rvalid = '1';
		wait for CLK_PERIOD_C;
		readDone_i           <= '0';
		counter_i            <= (others => '0');
		buffer_i             <= (others => (others => '0'));
		axiReadSrc_i.araddr  <= (others => '0');
		axiReadSrc_i.arlen   <= (others => '0');
		axiReadSrc_i.arsize  <= "000";
		axiReadSrc_i.arburst <= "00";
		axiReadSrc_i.arvalid <= '0';
		axiReadSrc_i.rready  <= '0';
		wait for CLK_PERIOD_C * 5;




		-- axi ready immediately, wait for data, read 2
		axiReadSrc_i.araddr  <= STD_LOGIC_VECTOR(to_unsigned(0, axiReadSrc_i.araddr'length));
		axiReadSrc_i.arlen   <= STD_LOGIC_VECTOR(to_unsigned(2-1, axiReadSrc_i.arlen'length));
		axiReadSrc_i.arsize  <= "101";
		axiReadSrc_i.arburst <= "01";
		axiReadSrc_i.arvalid <= '1';
		axiReadSrc_i.rready  <= '1';
		wait for CLK_PERIOD_C;
		axiReadSrc_i.arvalid <= '0';

		wait for CLK_PERIOD_C * 10;
		counter_i   <= to_unsigned(1, counter_i'length);
		buffer_i(0) <= x"badb17";
		wait for CLK_PERIOD_C;
		counter_i   <= to_unsigned(2, counter_i'length);
		buffer_i(1) <= x"ba5ad0";
		readDone_i  <= '1';

		--wait until axiReadDst_o.rvalid = '1';
		wait for CLK_PERIOD_C*2;
		readDone_i           <= '0';
		counter_i            <= (others => '0');
		buffer_i             <= (others => (others => '0'));
		axiReadSrc_i.araddr  <= (others => '0');
		axiReadSrc_i.arlen   <= (others => '0');
		axiReadSrc_i.arsize  <= "000";
		axiReadSrc_i.arburst <= "00";
		axiReadSrc_i.arvalid <= '0';
		axiReadSrc_i.rready  <= '0';
		wait for CLK_PERIOD_C * 5;




-- axi ready immediately, wait for data, read 3
		axiReadSrc_i.araddr  <= STD_LOGIC_VECTOR(to_unsigned(0, axiReadSrc_i.araddr'length));
		axiReadSrc_i.arlen   <= STD_LOGIC_VECTOR(to_unsigned(3-1, axiReadSrc_i.arlen'length));
		axiReadSrc_i.arsize  <= "101";
		axiReadSrc_i.arburst <= "01";
		axiReadSrc_i.arvalid <= '1';
		axiReadSrc_i.rready  <= '1';
		wait for CLK_PERIOD_C;
		axiReadSrc_i.arvalid <= '0';

		wait for CLK_PERIOD_C * 10;
		counter_i   <= to_unsigned(1, counter_i'length);
		buffer_i(0) <= x"badb17";
		wait for CLK_PERIOD_C;
		counter_i   <= to_unsigned(2, counter_i'length);
		buffer_i(1) <= x"baaaad";
		wait for CLK_PERIOD_C;
		counter_i   <= to_unsigned(3, counter_i'length);
		buffer_i(2) <= x"ba5ad0";
		readDone_i  <= '1';

		--wait until axiReadDst_o.rvalid = '1';
		wait for CLK_PERIOD_C*3;
		readDone_i           <= '0';
		counter_i            <= (others => '0');
		buffer_i             <= (others => (others => '0'));
		axiReadSrc_i.araddr  <= (others => '0');
		axiReadSrc_i.arlen   <= (others => '0');
		axiReadSrc_i.arsize  <= "000";
		axiReadSrc_i.arburst <= "00";
		axiReadSrc_i.arvalid <= '0';
		axiReadSrc_i.rready  <= '0';
		wait for CLK_PERIOD_C * 5;



		-- axi ready immediately, wait for data, read 4
		axiReadSrc_i.araddr  <= STD_LOGIC_VECTOR(to_unsigned(0, axiReadSrc_i.araddr'length));
		axiReadSrc_i.arlen   <= STD_LOGIC_VECTOR(to_unsigned(4-1, axiReadSrc_i.arlen'length));
		axiReadSrc_i.arsize  <= "101";
		axiReadSrc_i.arburst <= "01";
		axiReadSrc_i.arvalid <= '1';
		axiReadSrc_i.rready  <= '1';
		wait for CLK_PERIOD_C;
		axiReadSrc_i.arvalid <= '0';

		wait for CLK_PERIOD_C * 10;
		counter_i   <= to_unsigned(1, counter_i'length);
		buffer_i(0) <= x"badb17";
		wait for CLK_PERIOD_C;
		counter_i   <= to_unsigned(2, counter_i'length);
		buffer_i(1) <= x"baaaad";
		wait for CLK_PERIOD_C;
		counter_i   <= to_unsigned(3, counter_i'length);
		buffer_i(2) <= x"ba99ed";
		wait for CLK_PERIOD_C;
		counter_i   <= to_unsigned(0, counter_i'length);
		buffer_i(3) <= x"ba5ad0";
		readDone_i  <= '1';

		--wait until axiReadDst_o.rvalid = '1';
		wait for CLK_PERIOD_C*4;
		readDone_i           <= '0';
		counter_i            <= (others => '0');
		buffer_i             <= (others => (others => '0'));
		axiReadSrc_i.araddr  <= (others => '0');
		axiReadSrc_i.arlen   <= (others => '0');
		axiReadSrc_i.arsize  <= "000";
		axiReadSrc_i.arburst <= "00";
		axiReadSrc_i.arvalid <= '0';
		axiReadSrc_i.rready  <= '0';
		wait for CLK_PERIOD_C * 5;

		finish;

	end process stimulus;

end Behavioral;
